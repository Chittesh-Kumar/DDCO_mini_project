module tb_prefix_add8;
reg [7:0] t_a,t_b;
wire [7:0] t_sum;

prefix_add8 pa8 (.a(t_a), .b(t_b), .sum(t_sum));

initial begin $dumpfile("tb_prefix_add8.vcd"); 
$dumpvars(0, tb_prefix_add8); 
end

initial
begin
	t_a [7:0] = 8'b00000000; //0
	t_b [7:0] = 8'b01000001; //65
	
	#5
	t_a [7:0] = 8'b01100100; //100
	t_b [7:0] = 8'b00011000; //24

	#5
	t_a [7:0] = 8'b00010100; //20
	t_b [7:0] = 8'b10110010; //178
	
	#5
	t_a [7:0] = 8'b00100001; //33
	t_b [7:0] = 8'b00111111; //63
	
	#5
	t_a [7:0] = 8'b01100100; //100
	t_b [7:0] = 8'b00110010; //50
	
	#5
	t_a [7:0] = 8'b01100100; //100
	t_b [7:0] = 8'b00101000; //40

	#5
	t_a [7:0] = 8'b10110001; //177
	t_b [7:0] = 8'b00110110; //54
	
	#5
	t_a [7:0] = 8'b01011010; //90
	t_b [7:0] = 8'b00111100; //60
	
	#5
	t_a [7:0] = 8'b00011000; //24
	t_b [7:0] = 8'b01001100; //76
	
	#10
	t_a [7:0] = 8'b00000000;
	t_b [7:0] = 8'b00000001;
	#10
	t_a [7:0] = 8'b00000000;
	t_b [7:0] = 8'b00000001;
	
end
endmodule